module Rs();

endmodule;