module insCache(clk);
endmodule