module Rs();
endmodule;