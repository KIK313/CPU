module lsBuffer();
endmodule