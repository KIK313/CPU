module Rob(clk);
    input wire clk;
endmodule;