module ALU();
endmodule