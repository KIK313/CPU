module Rob();

endmodule;