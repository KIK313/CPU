module insFetch(
    input wire clk,
    input wire rst,
    input wire rdy,

    input wire[31:0] ins,
    output reg[31:0] ins_addr,
    
    
);


    always@ (posedge clk) begin
        if 
    end 

endmodule;