module insFetch(clk);
    input wire clk;
endmodule;