module memCtr (clk, rst, rdy, inData, outData);
    input wire clk;
    input wire rst;
    input wire rdy;
    input wire[7:0] inData;
    output reg[31:0] outData;
endmodule;