module regFile(clk);
    input wire clk;

endmodule