module Rs();

endmodule