module lsBuffer();
endmodule;